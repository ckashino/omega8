module cpu (clk, hold, opcode, d1, d2)
